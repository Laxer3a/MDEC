module GTEMicrocodeStart(
	input			IsNop,
	input	[5:0]	Instruction,
	output	[8:0]	StartAddress
);

	// TODO : Generate with C++ tool.

endmodule
