// Included file with constant : 
parameter
	// Bit 0 : Fist instruction -> Reset status bit.
	// Bit 1 : Last instruction -> Allow to end state.
	RSTFLG    = 59'b01,
	___FLG    = 59'b00,
	LAST__	  = 59'b10,
	
	// Bit 2 : Override and set to 0 the LM bit.
	USE_LM    = 1'b1,
	RST_LM    = 1'b0,
	// Bit  7:3
	// Bit 12:8
	DATA_VXY0 = 6'd0,
	DATA__VZ0 = 6'd1,
	DATA_VXY1 = 6'd2,
	DATA__VZ1 = 6'd3,
	DATA_VXY2 = 6'd4,
	DATA__VZ2 = 6'd5,
	DATA_RGBC = 6'd6,
	DATA__OTZ = 6'd7,
	DATA__IR0 = 6'd8,	D5TA_IR0 = 5'd8,
	DATA__IR1 = 6'd9,	D5TA_IR1 = 5'd9,
	DATA__IR2 = 6'd10,	D5TA_IR2 = 5'd10,
	DATA__IR3 = 6'd11,	D5TA_IR3 = 5'd11,
	DATA_SXY0 = 6'd12,
	DATA_SXY1 = 6'd13,
	DATA_SXY2 = 6'd14,
	DATA_SXYP = 6'd15,
	DATA__SZ0 = 6'd16,
	DATA__SZ1 = 6'd17,
	DATA__SZ2 = 6'd18,
	DATA__SZ3 = 6'd19,
	DATACRGB0 = 6'd20,
	DATACRGB1 = 6'd21,
	DATACRGB2 = 6'd22,
	DATA_RES1 = 6'd23,
	DATA_MAC0 = 6'd24,
	DATA_MAC1 = 6'd25,
	DATA_MAC2 = 6'd26,
	DATA_MAC3 = 6'd27,
	DATA_LZCR = 6'd30,
	
	DATA_STATUS = 5'd31,
	
	CT_R11R12 = 6'd32,
	CT_R13R21 = 6'd33,
	CT_R22R23 = 6'd34,
	CT_R31R32 = 6'd35,
	CT____R33 = 6'd36,
	CT_T_R_X_ = 6'd37,
	CT_T_R_Y_ = 6'd38,
	CT_T_R_Z_ = 6'd39,
	CT_L11L12 = 6'd40,
	CT_L13L21 = 6'd41,
	CT_L22L23 = 6'd42,
	CT_L31L32 = 6'd43,
	CT____L33 = 6'd44,
	CT_R_B_K_ = 6'd45,
	CT_G_B_K_ = 6'd46,
	CT_B_B_K_ = 6'd47,
	CT_LR1LR2 = 6'd48,
	CT_LR3LG1 = 6'd49,
	CT_LG2LG3 = 6'd50,
	CT_LB1LB2 = 6'd51,
	CT____LB3 = 6'd52,
	CT_R_F_C_ = 6'd53,
	CT_G_F_C_ = 6'd54,
	CT_B_F_C_ = 6'd55,
	CT_O_F_X_ = 6'd56,
	CT_O_F_Y_ = 6'd57,
	CT______H = 6'd58,
	CT____DQA = 6'd59,
	CT____DQB = 6'd60,
	CT___ZSF3 = 6'd61,
	CT___ZSF4 = 6'd62,
	
	DATA_____ = 6'd31,
	CTRL_____ = 6'd31,

	// WRITE
	DAT_WRITE = 1'b1,
	CTR_WRITE = 1'b1,
	____NOWRT = 1'b0,
	
	// Push
	PUSH___SZ = 1'b1,
	PUSH__SPX = 1'b1,
	PUSH__SPY = 1'b1,
	PUSH_CRGB = 1'b1,
	_NO_PSH__ = 1'b0,
	
	F______   = 19'b000_0000_0000_0000_0000,
	FLG_A1 	  = 19'b100_1000_0000_0000_0000,
	FLG_A2 	  = 19'b010_0100_0000_0000_0000,
	FLG_A3 	  = 19'b001_0010_0000_0000_0000,
	FLG_B1	  = 19'b000_0001_0000_0000_0000,
	FLG_B2	  = 19'b000_0000_1000_0000_0000,
	FLG_B3	  = 19'b000_0000_0100_0000_0000,
	
	UNUSED_SYMBOL_END_LIST = 0; // Convenience to add/remove item with the last , issue.
