// ----------------------------------------------------------------------------------------------
//   Compute Path
// ----------------------------------------------------------------------------------------------
`include "GTEDefine.hv"

module GTEComputePath(
	input					i_clk,
	input					i_nRst,
	
	input	CTRL			i_instrParam,
	input	gteComputeCtrl	i_computeCtrl,
	input	SgteREG			i_registers,
	output	gteCtrl			o_RegCtrl
);

	// [TODO Compute Path]

endmodule
