module InterpROM(
	input                clk,
	input         [ 8:0] adr,
	output signed [15:0] dataOut
);

reg [15:0] data;
assign dataOut = data;

always @(posedge clk) begin
	case (adr)
	9'd0  : data <= 16'hffff;
	9'd1  : data <= 16'hffff;
	9'd2  : data <= 16'hffff;
	9'd3  : data <= 16'hffff;
	9'd4  : data <= 16'hffff;
	9'd5  : data <= 16'hffff;
	9'd6  : data <= 16'hffff;
	9'd7  : data <= 16'hffff;
	9'd8  : data <= 16'hffff;
	9'd9  : data <= 16'hffff;
	9'd10 : data <= 16'hffff;
	9'd11 : data <= 16'hffff;
	9'd12 : data <= 16'hffff;
	9'd13 : data <= 16'hffff;
	9'd14 : data <= 16'hffff;
	9'd15 : data <= 16'hffff;
	9'd16 : data <= 16'h0;
	9'd17 : data <= 16'h0;
	9'd18 : data <= 16'h0;
	9'd19 : data <= 16'h0;
	9'd20 : data <= 16'h0;
	9'd21 : data <= 16'h0;
	9'd22 : data <= 16'h0;
	9'd23 : data <= 16'h1;
	9'd24 : data <= 16'h1;
	9'd25 : data <= 16'h1;
	9'd26 : data <= 16'h1;
	9'd27 : data <= 16'h2;
	9'd28 : data <= 16'h2;
	9'd29 : data <= 16'h2;
	9'd30 : data <= 16'h3;
	9'd31 : data <= 16'h3;
	9'd32 : data <= 16'h3;
	9'd33 : data <= 16'h4;
	9'd34 : data <= 16'h4;
	9'd35 : data <= 16'h5;
	9'd36 : data <= 16'h5;
	9'd37 : data <= 16'h6;
	9'd38 : data <= 16'h7;
	9'd39 : data <= 16'h7;
	9'd40 : data <= 16'h8;
	9'd41 : data <= 16'h9;
	9'd42 : data <= 16'h9;
	9'd43 : data <= 16'ha;
	9'd44 : data <= 16'hb;
	9'd45 : data <= 16'hc;
	9'd46 : data <= 16'hd;
	9'd47 : data <= 16'he;
	9'd48 : data <= 16'hf;
	9'd49 : data <= 16'h10;
	9'd50 : data <= 16'h11;
	9'd51 : data <= 16'h12;
	9'd52 : data <= 16'h13;
	9'd53 : data <= 16'h15;
	9'd54 : data <= 16'h16;
	9'd55 : data <= 16'h18;
	9'd56 : data <= 16'h19;
	9'd57 : data <= 16'h1b;
	9'd58 : data <= 16'h1c;
	9'd59 : data <= 16'h1e;
	9'd60 : data <= 16'h20;
	9'd61 : data <= 16'h21;
	9'd62 : data <= 16'h23;
	9'd63 : data <= 16'h25;
	9'd64 : data <= 16'h27;
	9'd65 : data <= 16'h29;
	9'd66 : data <= 16'h2c;
	9'd67 : data <= 16'h2e;
	9'd68 : data <= 16'h30;
	9'd69 : data <= 16'h33;
	9'd70 : data <= 16'h35;
	9'd71 : data <= 16'h38;
	9'd72 : data <= 16'h3a;
	9'd73 : data <= 16'h3d;
	9'd74 : data <= 16'h40;
	9'd75 : data <= 16'h43;
	9'd76 : data <= 16'h46;
	9'd77 : data <= 16'h49;
	9'd78 : data <= 16'h4d;
	9'd79 : data <= 16'h50;
	9'd80 : data <= 16'h54;
	9'd81 : data <= 16'h57;
	9'd82 : data <= 16'h5b;
	9'd83 : data <= 16'h5f;
	9'd84 : data <= 16'h63;
	9'd85 : data <= 16'h67;
	9'd86 : data <= 16'h6b;
	9'd87 : data <= 16'h6f;
	9'd88 : data <= 16'h74;
	9'd89 : data <= 16'h78;
	9'd90 : data <= 16'h7d;
	9'd91 : data <= 16'h82;
	9'd92 : data <= 16'h87;
	9'd93 : data <= 16'h8c;
	9'd94 : data <= 16'h91;
	9'd95 : data <= 16'h96;
	9'd96 : data <= 16'h9c;
	9'd97 : data <= 16'ha1;
	9'd98 : data <= 16'ha7;
	9'd99 : data <= 16'had;
	9'd100: data <= 16'hb3;
	9'd101: data <= 16'hba;
	9'd102: data <= 16'hc0;
	9'd103: data <= 16'hc7;
	9'd104: data <= 16'hcd;
	9'd105: data <= 16'hd4;
	9'd106: data <= 16'hdb;
	9'd107: data <= 16'he3;
	9'd108: data <= 16'hea;
	9'd109: data <= 16'hf2;
	9'd110: data <= 16'hfa;
	9'd111: data <= 16'h101;
	9'd112: data <= 16'h10a;
	9'd113: data <= 16'h112;
	9'd114: data <= 16'h11b;
	9'd115: data <= 16'h123;
	9'd116: data <= 16'h12c;
	9'd117: data <= 16'h135;
	9'd118: data <= 16'h13f;
	9'd119: data <= 16'h148;
	9'd120: data <= 16'h152;
	9'd121: data <= 16'h15c;
	9'd122: data <= 16'h166;
	9'd123: data <= 16'h171;
	9'd124: data <= 16'h17b;
	9'd125: data <= 16'h186;
	9'd126: data <= 16'h191;
	9'd127: data <= 16'h19c;
	9'd128: data <= 16'h1a8;
	9'd129: data <= 16'h1b4;
	9'd130: data <= 16'h1c0;
	9'd131: data <= 16'h1cc;
	9'd132: data <= 16'h1d9;
	9'd133: data <= 16'h1e5;
	9'd134: data <= 16'h1f2;
	9'd135: data <= 16'h200;
	9'd136: data <= 16'h20d;
	9'd137: data <= 16'h21b;
	9'd138: data <= 16'h229;
	9'd139: data <= 16'h237;
	9'd140: data <= 16'h246;
	9'd141: data <= 16'h255;
	9'd142: data <= 16'h264;
	9'd143: data <= 16'h273;
	9'd144: data <= 16'h283;
	9'd145: data <= 16'h293;
	9'd146: data <= 16'h2a3;
	9'd147: data <= 16'h2b4;
	9'd148: data <= 16'h2c4;
	9'd149: data <= 16'h2d6;
	9'd150: data <= 16'h2e7;
	9'd151: data <= 16'h2f9;
	9'd152: data <= 16'h30b;
	9'd153: data <= 16'h31d;
	9'd154: data <= 16'h330;
	9'd155: data <= 16'h343;
	9'd156: data <= 16'h356;
	9'd157: data <= 16'h36a;
	9'd158: data <= 16'h37e;
	9'd159: data <= 16'h392;
	9'd160: data <= 16'h3a7;
	9'd161: data <= 16'h3bc;
	9'd162: data <= 16'h3d1;
	9'd163: data <= 16'h3e7;
	9'd164: data <= 16'h3fc;
	9'd165: data <= 16'h413;
	9'd166: data <= 16'h42a;
	9'd167: data <= 16'h441;
	9'd168: data <= 16'h458;
	9'd169: data <= 16'h470;
	9'd170: data <= 16'h488;
	9'd171: data <= 16'h4a0;
	9'd172: data <= 16'h4b9;
	9'd173: data <= 16'h4d2;
	9'd174: data <= 16'h4ec;
	9'd175: data <= 16'h506;
	9'd176: data <= 16'h520;
	9'd177: data <= 16'h53b;
	9'd178: data <= 16'h556;
	9'd179: data <= 16'h572;
	9'd180: data <= 16'h58e;
	9'd181: data <= 16'h5aa;
	9'd182: data <= 16'h5c7;
	9'd183: data <= 16'h5e4;
	9'd184: data <= 16'h601;
	9'd185: data <= 16'h61f;
	9'd186: data <= 16'h63e;
	9'd187: data <= 16'h65c;
	9'd188: data <= 16'h67c;
	9'd189: data <= 16'h69b;
	9'd190: data <= 16'h6bb;
	9'd191: data <= 16'h6dc;
	9'd192: data <= 16'h6fd;
	9'd193: data <= 16'h71e;
	9'd194: data <= 16'h740;
	9'd195: data <= 16'h762;
	9'd196: data <= 16'h784;
	9'd197: data <= 16'h7a7;
	9'd198: data <= 16'h7cb;
	9'd199: data <= 16'h7ef;
	9'd200: data <= 16'h813;
	9'd201: data <= 16'h838;
	9'd202: data <= 16'h85d;
	9'd203: data <= 16'h883;
	9'd204: data <= 16'h8a9;
	9'd205: data <= 16'h8d0;
	9'd206: data <= 16'h8f7;
	9'd207: data <= 16'h91e;
	9'd208: data <= 16'h946;
	9'd209: data <= 16'h96f;
	9'd210: data <= 16'h998;
	9'd211: data <= 16'h9c1;
	9'd212: data <= 16'h9eb;
	9'd213: data <= 16'ha16;
	9'd214: data <= 16'ha40;
	9'd215: data <= 16'ha6c;
	9'd216: data <= 16'ha98;
	9'd217: data <= 16'hac4;
	9'd218: data <= 16'haf1;
	9'd219: data <= 16'hb1e;
	9'd220: data <= 16'hb4c;
	9'd221: data <= 16'hb7a;
	9'd222: data <= 16'hba9;
	9'd223: data <= 16'hbd8;
	9'd224: data <= 16'hc07;
	9'd225: data <= 16'hc38;
	9'd226: data <= 16'hc68;
	9'd227: data <= 16'hc99;
	9'd228: data <= 16'hccb;
	9'd229: data <= 16'hcfd;
	9'd230: data <= 16'hd30;
	9'd231: data <= 16'hd63;
	9'd232: data <= 16'hd97;
	9'd233: data <= 16'hdcb;
	9'd234: data <= 16'he00;
	9'd235: data <= 16'he35;
	9'd236: data <= 16'he6b;
	9'd237: data <= 16'hea1;
	9'd238: data <= 16'hed7;
	9'd239: data <= 16'hf0f;
	9'd240: data <= 16'hf46;
	9'd241: data <= 16'hf7f;
	9'd242: data <= 16'hfb7;
	9'd243: data <= 16'hff1;
	9'd244: data <= 16'h102a;
	9'd245: data <= 16'h1065;
	9'd246: data <= 16'h109f;
	9'd247: data <= 16'h10db;
	9'd248: data <= 16'h1116;
	9'd249: data <= 16'h1153;
	9'd250: data <= 16'h118f;
	9'd251: data <= 16'h11cd;
	9'd252: data <= 16'h120b;
	9'd253: data <= 16'h1249;
	9'd254: data <= 16'h1288;
	9'd255: data <= 16'h12c7;
	9'd256: data <= 16'h1307;
	9'd257: data <= 16'h1347;
	9'd258: data <= 16'h1388;
	9'd259: data <= 16'h13c9;
	9'd260: data <= 16'h140b;
	9'd261: data <= 16'h144d;
	9'd262: data <= 16'h1490;
	9'd263: data <= 16'h14d4;
	9'd264: data <= 16'h1517;
	9'd265: data <= 16'h155c;
	9'd266: data <= 16'h15a0;
	9'd267: data <= 16'h15e6;
	9'd268: data <= 16'h162c;
	9'd269: data <= 16'h1672;
	9'd270: data <= 16'h16b9;
	9'd271: data <= 16'h1700;
	9'd272: data <= 16'h1747;
	9'd273: data <= 16'h1790;
	9'd274: data <= 16'h17d8;
	9'd275: data <= 16'h1821;
	9'd276: data <= 16'h186b;
	9'd277: data <= 16'h18b5;
	9'd278: data <= 16'h1900;
	9'd279: data <= 16'h194b;
	9'd280: data <= 16'h1996;
	9'd281: data <= 16'h19e2;
	9'd282: data <= 16'h1a2e;
	9'd283: data <= 16'h1a7b;
	9'd284: data <= 16'h1ac8;
	9'd285: data <= 16'h1b16;
	9'd286: data <= 16'h1b64;
	9'd287: data <= 16'h1bb3;
	9'd288: data <= 16'h1c02;
	9'd289: data <= 16'h1c51;
	9'd290: data <= 16'h1ca1;
	9'd291: data <= 16'h1cf1;
	9'd292: data <= 16'h1d42;
	9'd293: data <= 16'h1d93;
	9'd294: data <= 16'h1de5;
	9'd295: data <= 16'h1e37;
	9'd296: data <= 16'h1e89;
	9'd297: data <= 16'h1edc;
	9'd298: data <= 16'h1f2f;
	9'd299: data <= 16'h1f82;
	9'd300: data <= 16'h1fd6;
	9'd301: data <= 16'h202a;
	9'd302: data <= 16'h207f;
	9'd303: data <= 16'h20d4;
	9'd304: data <= 16'h2129;
	9'd305: data <= 16'h217f;
	9'd306: data <= 16'h21d5;
	9'd307: data <= 16'h222c;
	9'd308: data <= 16'h2282;
	9'd309: data <= 16'h22da;
	9'd310: data <= 16'h2331;
	9'd311: data <= 16'h2389;
	9'd312: data <= 16'h23e1;
	9'd313: data <= 16'h2439;
	9'd314: data <= 16'h2492;
	9'd315: data <= 16'h24eb;
	9'd316: data <= 16'h2545;
	9'd317: data <= 16'h259e;
	9'd318: data <= 16'h25f8;
	9'd319: data <= 16'h2653;
	9'd320: data <= 16'h26ad;
	9'd321: data <= 16'h2708;
	9'd322: data <= 16'h2763;
	9'd323: data <= 16'h27be;
	9'd324: data <= 16'h281a;
	9'd325: data <= 16'h2876;
	9'd326: data <= 16'h28d2;
	9'd327: data <= 16'h292e;
	9'd328: data <= 16'h298b;
	9'd329: data <= 16'h29e7;
	9'd330: data <= 16'h2a44;
	9'd331: data <= 16'h2aa1;
	9'd332: data <= 16'h2aff;
	9'd333: data <= 16'h2b5c;
	9'd334: data <= 16'h2bba;
	9'd335: data <= 16'h2c18;
	9'd336: data <= 16'h2c76;
	9'd337: data <= 16'h2cd4;
	9'd338: data <= 16'h2d33;
	9'd339: data <= 16'h2d91;
	9'd340: data <= 16'h2df0;
	9'd341: data <= 16'h2e4f;
	9'd342: data <= 16'h2eae;
	9'd343: data <= 16'h2f0d;
	9'd344: data <= 16'h2f6c;
	9'd345: data <= 16'h2fcc;
	9'd346: data <= 16'h302b;
	9'd347: data <= 16'h308b;
	9'd348: data <= 16'h30ea;
	9'd349: data <= 16'h314a;
	9'd350: data <= 16'h31aa;
	9'd351: data <= 16'h3209;
	9'd352: data <= 16'h3269;
	9'd353: data <= 16'h32c9;
	9'd354: data <= 16'h3329;
	9'd355: data <= 16'h3389;
	9'd356: data <= 16'h33e9;
	9'd357: data <= 16'h3449;
	9'd358: data <= 16'h34a9;
	9'd359: data <= 16'h3509;
	9'd360: data <= 16'h3569;
	9'd361: data <= 16'h35c9;
	9'd362: data <= 16'h3629;
	9'd363: data <= 16'h3689;
	9'd364: data <= 16'h36e8;
	9'd365: data <= 16'h3748;
	9'd366: data <= 16'h37a8;
	9'd367: data <= 16'h3807;
	9'd368: data <= 16'h3867;
	9'd369: data <= 16'h38c6;
	9'd370: data <= 16'h3926;
	9'd371: data <= 16'h3985;
	9'd372: data <= 16'h39e4;
	9'd373: data <= 16'h3a43;
	9'd374: data <= 16'h3aa2;
	9'd375: data <= 16'h3b00;
	9'd376: data <= 16'h3b5f;
	9'd377: data <= 16'h3bbd;
	9'd378: data <= 16'h3c1b;
	9'd379: data <= 16'h3c79;
	9'd380: data <= 16'h3cd7;
	9'd381: data <= 16'h3d35;
	9'd382: data <= 16'h3d92;
	9'd383: data <= 16'h3def;
	9'd384: data <= 16'h3e4c;
	9'd385: data <= 16'h3ea9;
	9'd386: data <= 16'h3f05;
	9'd387: data <= 16'h3f62;
	9'd388: data <= 16'h3fbd;
	9'd389: data <= 16'h4019;
	9'd390: data <= 16'h4074;
	9'd391: data <= 16'h40d0;
	9'd392: data <= 16'h412a;
	9'd393: data <= 16'h4185;
	9'd394: data <= 16'h41df;
	9'd395: data <= 16'h4239;
	9'd396: data <= 16'h4292;
	9'd397: data <= 16'h42eb;
	9'd398: data <= 16'h4344;
	9'd399: data <= 16'h439c;
	9'd400: data <= 16'h43f4;
	9'd401: data <= 16'h444c;
	9'd402: data <= 16'h44a3;
	9'd403: data <= 16'h44fa;
	9'd404: data <= 16'h4550;
	9'd405: data <= 16'h45a6;
	9'd406: data <= 16'h45fc;
	9'd407: data <= 16'h4651;
	9'd408: data <= 16'h46a6;
	9'd409: data <= 16'h46fa;
	9'd410: data <= 16'h474e;
	9'd411: data <= 16'h47a1;
	9'd412: data <= 16'h47f4;
	9'd413: data <= 16'h4846;
	9'd414: data <= 16'h4898;
	9'd415: data <= 16'h48e9;
	9'd416: data <= 16'h493a;
	9'd417: data <= 16'h498a;
	9'd418: data <= 16'h49d9;
	9'd419: data <= 16'h4a29;
	9'd420: data <= 16'h4a77;
	9'd421: data <= 16'h4ac5;
	9'd422: data <= 16'h4b13;
	9'd423: data <= 16'h4b5f;
	9'd424: data <= 16'h4bac;
	9'd425: data <= 16'h4bf7;
	9'd426: data <= 16'h4c42;
	9'd427: data <= 16'h4c8d;
	9'd428: data <= 16'h4cd7;
	9'd429: data <= 16'h4d20;
	9'd430: data <= 16'h4d68;
	9'd431: data <= 16'h4db0;
	9'd432: data <= 16'h4df7;
	9'd433: data <= 16'h4e3e;
	9'd434: data <= 16'h4e84;
	9'd435: data <= 16'h4ec9;
	9'd436: data <= 16'h4f0e;
	9'd437: data <= 16'h4f52;
	9'd438: data <= 16'h4f95;
	9'd439: data <= 16'h4fd7;
	9'd440: data <= 16'h5019;
	9'd441: data <= 16'h505a;
	9'd442: data <= 16'h509a;
	9'd443: data <= 16'h50da;
	9'd444: data <= 16'h5118;
	9'd445: data <= 16'h5156;
	9'd446: data <= 16'h5194;
	9'd447: data <= 16'h51d0;
	9'd448: data <= 16'h520c;
	9'd449: data <= 16'h5247;
	9'd450: data <= 16'h5281;
	9'd451: data <= 16'h52ba;
	9'd452: data <= 16'h52f3;
	9'd453: data <= 16'h532a;
	9'd454: data <= 16'h5361;
	9'd455: data <= 16'h5397;
	9'd456: data <= 16'h53cc;
	9'd457: data <= 16'h5401;
	9'd458: data <= 16'h5434;
	9'd459: data <= 16'h5467;
	9'd460: data <= 16'h5499;
	9'd461: data <= 16'h54ca;
	9'd462: data <= 16'h54fa;
	9'd463: data <= 16'h5529;
	9'd464: data <= 16'h5558;
	9'd465: data <= 16'h5585;
	9'd466: data <= 16'h55b2;
	9'd467: data <= 16'h55de;
	9'd468: data <= 16'h5609;
	9'd469: data <= 16'h5632;
	9'd470: data <= 16'h565b;
	9'd471: data <= 16'h5684;
	9'd472: data <= 16'h56ab;
	9'd473: data <= 16'h56d1;
	9'd474: data <= 16'h56f6;
	9'd475: data <= 16'h571b;
	9'd476: data <= 16'h573e;
	9'd477: data <= 16'h5761;
	9'd478: data <= 16'h5782;
	9'd479: data <= 16'h57a3;
	9'd480: data <= 16'h57c3;
	9'd481: data <= 16'h57e2;
	9'd482: data <= 16'h57ff;
	9'd483: data <= 16'h581c;
	9'd484: data <= 16'h5838;
	9'd485: data <= 16'h5853;
	9'd486: data <= 16'h586d;
	9'd487: data <= 16'h5886;
	9'd488: data <= 16'h589e;
	9'd489: data <= 16'h58b5;
	9'd490: data <= 16'h58cb;
	9'd491: data <= 16'h58e0;
	9'd492: data <= 16'h58f4;
	9'd493: data <= 16'h5907;
	9'd494: data <= 16'h5919;
	9'd495: data <= 16'h592a;
	9'd496: data <= 16'h593a;
	9'd497: data <= 16'h5949;
	9'd498: data <= 16'h5958;
	9'd499: data <= 16'h5965;
	9'd500: data <= 16'h5971;
	9'd501: data <= 16'h597c;
	9'd502: data <= 16'h5986;
	9'd503: data <= 16'h598f;
	9'd504: data <= 16'h5997;
	9'd505: data <= 16'h599e;
	9'd506: data <= 16'h59a4;
	9'd507: data <= 16'h59a9;
	9'd508: data <= 16'h59ad;
	9'd509: data <= 16'h59b0;
	9'd510: data <= 16'h59b2;
	9'd511: data <= 16'h59b3;
	endcase
end
	
endmodule
