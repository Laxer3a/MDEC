// ----------------------------------------------------------------------------------------------
//   Microcode RAM/ROM
// ----------------------------------------------------------------------------------------------
`include "GTEDefine.hv"

module GTEMicroCode(
	input					i_clk,
	input [8:0]				i_PC,
	
	output gteComputeCtrl	o_ctrl,
	output o_lastInstr
);

	// [TODO Microcode Generator]

endmodule
