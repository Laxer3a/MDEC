module FileReg (
	input         clk,
	input         read,
	input   [4:0] readAdr,
	output [31:0] outData,
	input         write,
	input   [4:0] writeAdr,
	input  [31:0] inData
);

	// TODO
	
endmodule